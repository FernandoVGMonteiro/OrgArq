library ieee;
use ieee.std_logic_1164.ALL;
use ieee.numeric_std.all;

entity instruction_cache is
port (clock: in std_logic;
		address: in  std_logic_vector(31 downto 0);
		dataOut: out std_logic_vector(31 downto 0)
		);
end entity;

architecture arch of instruction_cache is

type cache_data is array (0 to 15) of std_logic_vector(31 downto 0);
constant cache: cache_data := (
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000"
	);

signal addressInt: integer;
	
begin
	
	addressInt <= to_integer(unsigned(address));
	dataOut <= cache(addressInt);

end architecture;